`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////
// Institution:    Universidade Federal de Sergipe
// Engineer:       Saulo G. Felix
//
// Create Date:    02:54:35 09/30/2019
// Design Name:    Saulo G. Felix
// Module Name:    fifo_memory_unit
// Project Name:   elevetor_controller
// Target Devices: Spartan3E
// Tool versions:  ISE 14.7
// Description:    FIFO Memory queue
///////////////////////////////////////////////////////////////////////////////
module fifo_memory_unit(
    );

endmodule
