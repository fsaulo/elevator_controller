`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:        Universidade Federal de Sergipe
// Engineer:       
// 
// Create Date:    10:22:52 09/26/2019 
// Design Name:    Saulo G. Felix
// Module Name:    control_input_module 
// Project Name:   elevetor_controller
// Target Devices: Spartan3E
// Tool versions:  ISE 14.7
// Description:    The control system module
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module control_input_module(
    );


endmodule
